** Profile: "SCHEMATIC1-test"  [ E:\Tehnici CAD\proiect\proiectcad_sabauradubogdan-pspicefiles\schematic1\test.sim ] 

** Creating circuit file "test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ledorange.lib" 
* From [PSPICE NETLIST] section of E:\CAD\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.MC 5 TRAN V([OUT]) YMAX OUTPUT ALL SEED=200 
.STEP LIN PARAM R 22k 32k 2k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
